-- Javier Otero Martinez
-- OctaveSax project -- TFG
-- June 2019

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity istft_window_rom is Port (
	in_frame : in STD_LOGIC_VECTOR(8 downto 0);
	out_win : out STD_LOGIC_VECTOR(15 downto 0)
	);
end istft_window_rom;

architecture Behavioral of istft_window_rom is

	begin

	with in_frame select out_win <=
		"0000000000000000" when "000000001",
		"0000000000000011" when "000000010",
		"0000000000000111" when "000000011",
		"0000000000001101" when "000000100",
		"0000000000010100" when "000000101",
		"0000000000011101" when "000000110",
		"0000000000101000" when "000000111",
		"0000000000110100" when "000001000",
		"0000000001000010" when "000001001",
		"0000000001010010" when "000001010",
		"0000000001100011" when "000001011",
		"0000000001110110" when "000001100",
		"0000000010001010" when "000001101",
		"0000000010100000" when "000001110",
		"0000000010111000" when "000001111",
		"0000000011010001" when "000010000",
		"0000000011101100" when "000010001",
		"0000000100001001" when "000010010",
		"0000000100100111" when "000010011",
		"0000000101000111" when "000010100",
		"0000000101101000" when "000010101",
		"0000000110001011" when "000010110",
		"0000000110110000" when "000010111",
		"0000000111010110" when "000011000",
		"0000000111111110" when "000011001",
		"0000001000100111" when "000011010",
		"0000001001010010" when "000011011",
		"0000001001111110" when "000011100",
		"0000001010101100" when "000011101",
		"0000001011011011" when "000011110",
		"0000001100001100" when "000011111",
		"0000001100111111" when "000100000",
		"0000001101110011" when "000100001",
		"0000001110101001" when "000100010",
		"0000001111100000" when "000100011",
		"0000010000011000" when "000100100",
		"0000010001010010" when "000100101",
		"0000010010001110" when "000100110",
		"0000010011001011" when "000100111",
		"0000010100001001" when "000101000",
		"0000010101001001" when "000101001",
		"0000010110001010" when "000101010",
		"0000010111001101" when "000101011",
		"0000011000010001" when "000101100",
		"0000011001010111" when "000101101",
		"0000011010011110" when "000101110",
		"0000011011100111" when "000101111",
		"0000011100110000" when "000110000",
		"0000011101111011" when "000110001",
		"0000011111001000" when "000110010",
		"0000100000010110" when "000110011",
		"0000100001100101" when "000110100",
		"0000100010110110" when "000110101",
		"0000100100000111" when "000110110",
		"0000100101011010" when "000110111",
		"0000100110101111" when "000111000",
		"0000101000000100" when "000111001",
		"0000101001011011" when "000111010",
		"0000101010110100" when "000111011",
		"0000101100001101" when "000111100",
		"0000101101101000" when "000111101",
		"0000101111000011" when "000111110",
		"0000110000100000" when "000111111",
		"0000110001111111" when "001000000",
		"0000110011011110" when "001000001",
		"0000110100111111" when "001000010",
		"0000110110100000" when "001000011",
		"0000111000000011" when "001000100",
		"0000111001100111" when "001000101",
		"0000111011001100" when "001000110",
		"0000111100110010" when "001000111",
		"0000111110011001" when "001001000",
		"0001000000000001" when "001001001",
		"0001000001101010" when "001001010",
		"0001000011010100" when "001001011",
		"0001000101000000" when "001001100",
		"0001000110101100" when "001001101",
		"0001001000011001" when "001001110",
		"0001001010000111" when "001001111",
		"0001001011110110" when "001010000",
		"0001001101100110" when "001010001",
		"0001001111010111" when "001010010",
		"0001010001001000" when "001010011",
		"0001010010111011" when "001010100",
		"0001010100101110" when "001010101",
		"0001010110100010" when "001010110",
		"0001011000010111" when "001010111",
		"0001011010001101" when "001011000",
		"0001011100000100" when "001011001",
		"0001011101111011" when "001011010",
		"0001011111110011" when "001011011",
		"0001100001101100" when "001011100",
		"0001100011100110" when "001011101",
		"0001100101100000" when "001011110",
		"0001100111011011" when "001011111",
		"0001101001010110" when "001100000",
		"0001101011010010" when "001100001",
		"0001101101001111" when "001100010",
		"0001101111001101" when "001100011",
		"0001110001001010" when "001100100",
		"0001110011001001" when "001100101",
		"0001110101001000" when "001100110",
		"0001110111000111" when "001100111",
		"0001111001000111" when "001101000",
		"0001111011001000" when "001101001",
		"0001111101001001" when "001101010",
		"0001111111001010" when "001101011",
		"0010000001001100" when "001101100",
		"0010000011001110" when "001101101",
		"0010000101010001" when "001101110",
		"0010000111010100" when "001101111",
		"0010001001010111" when "001110000",
		"0010001011011011" when "001110001",
		"0010001101011111" when "001110010",
		"0010001111100011" when "001110011",
		"0010010001100111" when "001110100",
		"0010010011101100" when "001110101",
		"0010010101110001" when "001110110",
		"0010010111110110" when "001110111",
		"0010011001111100" when "001111000",
		"0010011100000001" when "001111001",
		"0010011110000111" when "001111010",
		"0010100000001100" when "001111011",
		"0010100010010010" when "001111100",
		"0010100100011000" when "001111101",
		"0010100110011110" when "001111110",
		"0010101000100100" when "001111111",
		"0010101010101010" when "010000000",
		"0010101100110000" when "010000001",
		"0010101110110110" when "010000010",
		"0010110000111100" when "010000011",
		"0010110011000010" when "010000100",
		"0010110101001000" when "010000101",
		"0010110111001110" when "010000110",
		"0010111001010011" when "010000111",
		"0010111011011001" when "010001000",
		"0010111101011110" when "010001001",
		"0010111111100011" when "010001010",
		"0011000001101000" when "010001011",
		"0011000011101101" when "010001100",
		"0011000101110001" when "010001101",
		"0011000111110110" when "010001110",
		"0011001001111001" when "010001111",
		"0011001011111101" when "010010000",
		"0011001110000000" when "010010001",
		"0011010000000011" when "010010010",
		"0011010010000110" when "010010011",
		"0011010100001000" when "010010100",
		"0011010110001010" when "010010101",
		"0011011000001011" when "010010110",
		"0011011010001100" when "010010111",
		"0011011100001101" when "010011000",
		"0011011110001101" when "010011001",
		"0011100000001100" when "010011010",
		"0011100010001011" when "010011011",
		"0011100100001010" when "010011100",
		"0011100110001000" when "010011101",
		"0011101000000101" when "010011110",
		"0011101010000010" when "010011111",
		"0011101011111110" when "010100000",
		"0011101101111010" when "010100001",
		"0011101111110100" when "010100010",
		"0011110001101111" when "010100011",
		"0011110011101000" when "010100100",
		"0011110101100001" when "010100101",
		"0011110111011001" when "010100110",
		"0011111001010000" when "010100111",
		"0011111011000111" when "010101000",
		"0011111100111101" when "010101001",
		"0011111110110010" when "010101010",
		"0100000000100110" when "010101011",
		"0100000010011010" when "010101100",
		"0100000100001100" when "010101101",
		"0100000101111110" when "010101110",
		"0100000111101111" when "010101111",
		"0100001001011110" when "010110000",
		"0100001011001101" when "010110001",
		"0100001100111100" when "010110010",
		"0100001110101001" when "010110011",
		"0100010000010101" when "010110100",
		"0100010010000000" when "010110101",
		"0100010011101010" when "010110110",
		"0100010101010011" when "010110111",
		"0100010110111011" when "010111000",
		"0100011000100011" when "010111001",
		"0100011010001001" when "010111010",
		"0100011011101110" when "010111011",
		"0100011101010001" when "010111100",
		"0100011110110100" when "010111101",
		"0100100000010110" when "010111110",
		"0100100001110110" when "010111111",
		"0100100011010110" when "011000000",
		"0100100100110100" when "011000001",
		"0100100110010001" when "011000010",
		"0100100111101101" when "011000011",
		"0100101001000111" when "011000100",
		"0100101010100001" when "011000101",
		"0100101011111001" when "011000110",
		"0100101101010000" when "011000111",
		"0100101110100110" when "011001000",
		"0100101111111010" when "011001001",
		"0100110001001101" when "011001010",
		"0100110010011111" when "011001011",
		"0100110011101111" when "011001100",
		"0100110100111111" when "011001101",
		"0100110110001100" when "011001110",
		"0100110111011001" when "011001111",
		"0100111000100100" when "011010000",
		"0100111001101110" when "011010001",
		"0100111010110110" when "011010010",
		"0100111011111101" when "011010011",
		"0100111101000011" when "011010100",
		"0100111110000111" when "011010101",
		"0100111111001010" when "011010110",
		"0101000000001011" when "011010111",
		"0101000001001011" when "011011000",
		"0101000010001010" when "011011001",
		"0101000011000111" when "011011010",
		"0101000100000010" when "011011011",
		"0101000100111100" when "011011100",
		"0101000101110101" when "011011101",
		"0101000110101100" when "011011110",
		"0101000111100001" when "011011111",
		"0101001000010101" when "011100000",
		"0101001001001000" when "011100001",
		"0101001001111001" when "011100010",
		"0101001010101000" when "011100011",
		"0101001011010110" when "011100100",
		"0101001100000011" when "011100101",
		"0101001100101110" when "011100110",
		"0101001101010111" when "011100111",
		"0101001101111111" when "011101000",
		"0101001110100101" when "011101001",
		"0101001111001001" when "011101010",
		"0101001111101100" when "011101011",
		"0101010000001101" when "011101100",
		"0101010000101101" when "011101101",
		"0101010001001011" when "011101110",
		"0101010001101000" when "011101111",
		"0101010010000011" when "011110000",
		"0101010010011100" when "011110001",
		"0101010010110100" when "011110010",
		"0101010011001010" when "011110011",
		"0101010011011111" when "011110100",
		"0101010011110001" when "011110101",
		"0101010100000011" when "011110110",
		"0101010100010010" when "011110111",
		"0101010100100000" when "011111000",
		"0101010100101101" when "011111001",
		"0101010100110111" when "011111010",
		"0101010101000000" when "011111011",
		"0101010101001000" when "011111100",
		"0101010101001101" when "011111101",
		"0101010101010010" when "011111110",
		"0101010101010100" when "011111111",
		"0101010101010101" when "100000000",
		"0101010101010100" when "100000001",
		"0101010101010010" when "100000010",
		"0101010101001101" when "100000011",
		"0101010101001000" when "100000100",
		"0101010101000000" when "100000101",
		"0101010100110111" when "100000110",
		"0101010100101101" when "100000111",
		"0101010100100000" when "100001000",
		"0101010100010010" when "100001001",
		"0101010100000011" when "100001010",
		"0101010011110001" when "100001011",
		"0101010011011111" when "100001100",
		"0101010011001010" when "100001101",
		"0101010010110100" when "100001110",
		"0101010010011100" when "100001111",
		"0101010010000011" when "100010000",
		"0101010001101000" when "100010001",
		"0101010001001011" when "100010010",
		"0101010000101101" when "100010011",
		"0101010000001101" when "100010100",
		"0101001111101100" when "100010101",
		"0101001111001001" when "100010110",
		"0101001110100101" when "100010111",
		"0101001101111111" when "100011000",
		"0101001101010111" when "100011001",
		"0101001100101110" when "100011010",
		"0101001100000011" when "100011011",
		"0101001011010110" when "100011100",
		"0101001010101000" when "100011101",
		"0101001001111001" when "100011110",
		"0101001001001000" when "100011111",
		"0101001000010101" when "100100000",
		"0101000111100001" when "100100001",
		"0101000110101100" when "100100010",
		"0101000101110101" when "100100011",
		"0101000100111100" when "100100100",
		"0101000100000010" when "100100101",
		"0101000011000111" when "100100110",
		"0101000010001010" when "100100111",
		"0101000001001011" when "100101000",
		"0101000000001011" when "100101001",
		"0100111111001010" when "100101010",
		"0100111110000111" when "100101011",
		"0100111101000011" when "100101100",
		"0100111011111101" when "100101101",
		"0100111010110110" when "100101110",
		"0100111001101110" when "100101111",
		"0100111000100100" when "100110000",
		"0100110111011001" when "100110001",
		"0100110110001100" when "100110010",
		"0100110100111111" when "100110011",
		"0100110011101111" when "100110100",
		"0100110010011111" when "100110101",
		"0100110001001101" when "100110110",
		"0100101111111010" when "100110111",
		"0100101110100110" when "100111000",
		"0100101101010000" when "100111001",
		"0100101011111001" when "100111010",
		"0100101010100001" when "100111011",
		"0100101001000111" when "100111100",
		"0100100111101101" when "100111101",
		"0100100110010001" when "100111110",
		"0100100100110100" when "100111111",
		"0100100011010110" when "101000000",
		"0100100001110110" when "101000001",
		"0100100000010110" when "101000010",
		"0100011110110100" when "101000011",
		"0100011101010001" when "101000100",
		"0100011011101110" when "101000101",
		"0100011010001001" when "101000110",
		"0100011000100011" when "101000111",
		"0100010110111011" when "101001000",
		"0100010101010011" when "101001001",
		"0100010011101010" when "101001010",
		"0100010010000000" when "101001011",
		"0100010000010101" when "101001100",
		"0100001110101001" when "101001101",
		"0100001100111100" when "101001110",
		"0100001011001101" when "101001111",
		"0100001001011110" when "101010000",
		"0100000111101111" when "101010001",
		"0100000101111110" when "101010010",
		"0100000100001100" when "101010011",
		"0100000010011010" when "101010100",
		"0100000000100110" when "101010101",
		"0011111110110010" when "101010110",
		"0011111100111101" when "101010111",
		"0011111011000111" when "101011000",
		"0011111001010000" when "101011001",
		"0011110111011001" when "101011010",
		"0011110101100001" when "101011011",
		"0011110011101000" when "101011100",
		"0011110001101111" when "101011101",
		"0011101111110100" when "101011110",
		"0011101101111010" when "101011111",
		"0011101011111110" when "101100000",
		"0011101010000010" when "101100001",
		"0011101000000101" when "101100010",
		"0011100110001000" when "101100011",
		"0011100100001010" when "101100100",
		"0011100010001011" when "101100101",
		"0011100000001100" when "101100110",
		"0011011110001101" when "101100111",
		"0011011100001101" when "101101000",
		"0011011010001100" when "101101001",
		"0011011000001011" when "101101010",
		"0011010110001010" when "101101011",
		"0011010100001000" when "101101100",
		"0011010010000110" when "101101101",
		"0011010000000011" when "101101110",
		"0011001110000000" when "101101111",
		"0011001011111101" when "101110000",
		"0011001001111001" when "101110001",
		"0011000111110110" when "101110010",
		"0011000101110001" when "101110011",
		"0011000011101101" when "101110100",
		"0011000001101000" when "101110101",
		"0010111111100011" when "101110110",
		"0010111101011110" when "101110111",
		"0010111011011001" when "101111000",
		"0010111001010011" when "101111001",
		"0010110111001110" when "101111010",
		"0010110101001000" when "101111011",
		"0010110011000010" when "101111100",
		"0010110000111100" when "101111101",
		"0010101110110110" when "101111110",
		"0010101100110000" when "101111111",
		"0010101010101010" when "110000000",
		"0010101000100100" when "110000001",
		"0010100110011110" when "110000010",
		"0010100100011000" when "110000011",
		"0010100010010010" when "110000100",
		"0010100000001100" when "110000101",
		"0010011110000111" when "110000110",
		"0010011100000001" when "110000111",
		"0010011001111100" when "110001000",
		"0010010111110110" when "110001001",
		"0010010101110001" when "110001010",
		"0010010011101100" when "110001011",
		"0010010001100111" when "110001100",
		"0010001111100011" when "110001101",
		"0010001101011111" when "110001110",
		"0010001011011011" when "110001111",
		"0010001001010111" when "110010000",
		"0010000111010100" when "110010001",
		"0010000101010001" when "110010010",
		"0010000011001110" when "110010011",
		"0010000001001100" when "110010100",
		"0001111111001010" when "110010101",
		"0001111101001001" when "110010110",
		"0001111011001000" when "110010111",
		"0001111001000111" when "110011000",
		"0001110111000111" when "110011001",
		"0001110101001000" when "110011010",
		"0001110011001001" when "110011011",
		"0001110001001010" when "110011100",
		"0001101111001101" when "110011101",
		"0001101101001111" when "110011110",
		"0001101011010010" when "110011111",
		"0001101001010110" when "110100000",
		"0001100111011011" when "110100001",
		"0001100101100000" when "110100010",
		"0001100011100110" when "110100011",
		"0001100001101100" when "110100100",
		"0001011111110011" when "110100101",
		"0001011101111011" when "110100110",
		"0001011100000100" when "110100111",
		"0001011010001101" when "110101000",
		"0001011000010111" when "110101001",
		"0001010110100010" when "110101010",
		"0001010100101110" when "110101011",
		"0001010010111011" when "110101100",
		"0001010001001000" when "110101101",
		"0001001111010111" when "110101110",
		"0001001101100110" when "110101111",
		"0001001011110110" when "110110000",
		"0001001010000111" when "110110001",
		"0001001000011001" when "110110010",
		"0001000110101100" when "110110011",
		"0001000101000000" when "110110100",
		"0001000011010100" when "110110101",
		"0001000001101010" when "110110110",
		"0001000000000001" when "110110111",
		"0000111110011001" when "110111000",
		"0000111100110010" when "110111001",
		"0000111011001100" when "110111010",
		"0000111001100111" when "110111011",
		"0000111000000011" when "110111100",
		"0000110110100000" when "110111101",
		"0000110100111111" when "110111110",
		"0000110011011110" when "110111111",
		"0000110001111111" when "111000000",
		"0000110000100000" when "111000001",
		"0000101111000011" when "111000010",
		"0000101101101000" when "111000011",
		"0000101100001101" when "111000100",
		"0000101010110100" when "111000101",
		"0000101001011011" when "111000110",
		"0000101000000100" when "111000111",
		"0000100110101111" when "111001000",
		"0000100101011010" when "111001001",
		"0000100100000111" when "111001010",
		"0000100010110110" when "111001011",
		"0000100001100101" when "111001100",
		"0000100000010110" when "111001101",
		"0000011111001000" when "111001110",
		"0000011101111011" when "111001111",
		"0000011100110000" when "111010000",
		"0000011011100111" when "111010001",
		"0000011010011110" when "111010010",
		"0000011001010111" when "111010011",
		"0000011000010001" when "111010100",
		"0000010111001101" when "111010101",
		"0000010110001010" when "111010110",
		"0000010101001001" when "111010111",
		"0000010100001001" when "111011000",
		"0000010011001011" when "111011001",
		"0000010010001110" when "111011010",
		"0000010001010010" when "111011011",
		"0000010000011000" when "111011100",
		"0000001111100000" when "111011101",
		"0000001110101001" when "111011110",
		"0000001101110011" when "111011111",
		"0000001100111111" when "111100000",
		"0000001100001100" when "111100001",
		"0000001011011011" when "111100010",
		"0000001010101100" when "111100011",
		"0000001001111110" when "111100100",
		"0000001001010010" when "111100101",
		"0000001000100111" when "111100110",
		"0000000111111110" when "111100111",
		"0000000111010110" when "111101000",
		"0000000110110000" when "111101001",
		"0000000110001011" when "111101010",
		"0000000101101000" when "111101011",
		"0000000101000111" when "111101100",
		"0000000100100111" when "111101101",
		"0000000100001001" when "111101110",
		"0000000011101100" when "111101111",
		"0000000011010001" when "111110000",
		"0000000010111000" when "111110001",
		"0000000010100000" when "111110010",
		"0000000010001010" when "111110011",
		"0000000001110110" when "111110100",
		"0000000001100011" when "111110101",
		"0000000001010010" when "111110110",
		"0000000001000010" when "111110111",
		"0000000000110100" when "111111000",
		"0000000000101000" when "111111001",
		"0000000000011101" when "111111010",
		"0000000000010100" when "111111011",
		"0000000000001101" when "111111100",
		"0000000000000111" when "111111101",
		"0000000000000011" when "111111110",
		"0000000000000000" when "111111111",
		"0000000000000000" when others;
end Behavioral